module spi()

endmodule